//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Top-level Verilog module for FPGA
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Fri Sep  5 11:54:22 2025
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
`default_nettype none

// ----- Verilog module for fpga_top -----
module fpga_top(pReset,
                prog_clk,
                set,
                reset,
                clk,
                gfpga_pad_GPIO_PAD,
                ccff_head,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] pReset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- GLOBAL PORTS -----
input [0:0] set;
//----- GLOBAL PORTS -----
input [0:0] reset;
//----- GLOBAL PORTS -----
input [0:0] clk;
//----- GPIO PORTS -----
inout [0:63] gfpga_pad_GPIO_PAD;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__0_ccff_tail;
wire [0:10] cbx_1__0__0_chanx_left_out;
wire [0:10] cbx_1__0__0_chanx_right_out;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_1__1__0_ccff_tail;
wire [0:10] cbx_1__1__0_chanx_left_out;
wire [0:10] cbx_1__1__0_chanx_right_out;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_;
wire [0:0] cbx_1__2__0_ccff_tail;
wire [0:10] cbx_1__2__0_chanx_left_out;
wire [0:10] cbx_1__2__0_chanx_right_out;
wire [0:0] cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__2__1_ccff_tail;
wire [0:10] cbx_1__2__1_chanx_left_out;
wire [0:10] cbx_1__2__1_chanx_right_out;
wire [0:0] cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_2__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_2__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_2__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_2__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_2__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_2__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_2__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_2__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_2__0__0_ccff_tail;
wire [0:10] cbx_2__0__0_chanx_left_out;
wire [0:10] cbx_2__0__0_chanx_right_out;
wire [0:0] cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_4_;
wire [0:0] cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_5_;
wire [0:0] cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_6_;
wire [0:0] cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_7_;
wire [0:0] cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_5_;
wire [0:0] cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_6_;
wire [0:0] cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_7_;
wire [0:0] cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_8_;
wire [0:0] cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_9_;
wire [0:0] cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ren_0_;
wire [0:0] cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_5_;
wire [0:0] cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_6_;
wire [0:0] cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_7_;
wire [0:0] cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_8_;
wire [0:0] cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_9_;
wire [0:0] cby_0__1__0_ccff_tail;
wire [0:10] cby_0__1__0_chany_bottom_out;
wire [0:10] cby_0__1__0_chany_top_out;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] cby_0__1__1_ccff_tail;
wire [0:10] cby_0__1__1_chany_bottom_out;
wire [0:10] cby_0__1__1_chany_top_out;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] cby_1__1__0_ccff_tail;
wire [0:10] cby_1__1__0_chany_bottom_out;
wire [0:10] cby_1__1__0_chany_top_out;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] cby_1__2__0_ccff_tail;
wire [0:10] cby_1__2__0_chany_bottom_out;
wire [0:10] cby_1__2__0_chany_top_out;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_18_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_19_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_2__1__0_ccff_tail;
wire [0:10] cby_2__1__0_chany_bottom_out;
wire [0:10] cby_2__1__0_chany_top_out;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_data_in_1_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_data_in_2_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_data_in_3_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_raddr_0_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_raddr_2_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_raddr_3_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_raddr_4_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_waddr_0_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_waddr_1_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_waddr_3_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_waddr_4_;
wire [0:0] cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_;
wire [0:0] cby_2__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_2__1__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_2__1__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_2__1__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_2__1__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_2__1__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_2__1__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_2__1__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_2__2__0_ccff_tail;
wire [0:10] cby_2__2__0_chany_bottom_out;
wire [0:10] cby_2__2__0_chany_top_out;
wire [0:0] cby_2__2__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_2__2__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_2__2__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_2__2__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_2__2__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_2__2__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_2__2__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_2__2__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_0_ccff_tail;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_1__1__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_;
wire [0:0] grid_clb_1__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_10_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_11_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_12_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_13_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_14_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_15_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_16_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_17_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_18_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_19_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_4_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_5_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_6_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_7_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_;
wire [0:0] grid_io_bottom_0_ccff_tail;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_ccff_tail;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_0_ccff_tail;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_1_ccff_tail;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_0_ccff_tail;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_1_ccff_tail;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_0_ccff_tail;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_1_ccff_tail;
wire [0:0] grid_memory_0_bottom_width_0_height_0_subtile_0__pin_data_out_4_;
wire [0:0] grid_memory_0_bottom_width_0_height_0_subtile_0__pin_data_out_5_;
wire [0:0] grid_memory_0_bottom_width_0_height_0_subtile_0__pin_data_out_6_;
wire [0:0] grid_memory_0_bottom_width_0_height_0_subtile_0__pin_data_out_7_;
wire [0:0] grid_memory_0_right_width_0_height_0_subtile_0__pin_data_out_0_;
wire [0:0] grid_memory_0_right_width_0_height_0_subtile_0__pin_data_out_1_;
wire [0:0] grid_memory_0_right_width_0_height_0_subtile_0__pin_data_out_2_;
wire [0:0] grid_memory_0_right_width_0_height_0_subtile_0__pin_data_out_3_;
wire [0:0] sb_0__0__0_ccff_tail;
wire [0:10] sb_0__0__0_chanx_right_out;
wire [0:10] sb_0__0__0_chany_top_out;
wire [0:0] sb_0__1__0_ccff_tail;
wire [0:10] sb_0__1__0_chanx_right_out;
wire [0:10] sb_0__1__0_chany_bottom_out;
wire [0:10] sb_0__1__0_chany_top_out;
wire [0:0] sb_0__2__0_ccff_tail;
wire [0:10] sb_0__2__0_chanx_right_out;
wire [0:10] sb_0__2__0_chany_bottom_out;
wire [0:0] sb_1__0__0_ccff_tail;
wire [0:10] sb_1__0__0_chanx_left_out;
wire [0:10] sb_1__0__0_chanx_right_out;
wire [0:10] sb_1__0__0_chany_top_out;
wire [0:0] sb_1__1__0_ccff_tail;
wire [0:10] sb_1__1__0_chanx_left_out;
wire [0:10] sb_1__1__0_chany_bottom_out;
wire [0:10] sb_1__1__0_chany_top_out;
wire [0:0] sb_1__2__0_ccff_tail;
wire [0:10] sb_1__2__0_chanx_left_out;
wire [0:10] sb_1__2__0_chanx_right_out;
wire [0:10] sb_1__2__0_chany_bottom_out;
wire [0:0] sb_2__0__0_ccff_tail;
wire [0:10] sb_2__0__0_chanx_left_out;
wire [0:10] sb_2__0__0_chany_top_out;
wire [0:0] sb_2__1__0_ccff_tail;
wire [0:10] sb_2__1__0_chany_bottom_out;
wire [0:10] sb_2__1__0_chany_top_out;
wire [0:0] sb_2__2__0_ccff_tail;
wire [0:10] sb_2__2__0_chanx_left_out;
wire [0:10] sb_2__2__0_chany_bottom_out;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	grid_io_top grid_io_top_1__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[0:7]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__2__0_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_0_ccff_tail));

	grid_io_top grid_io_top_2__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[8:15]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__2__1_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_1_ccff_tail));

	grid_io_right grid_io_right_3__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[16:23]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_2__2__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_2__2__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_2__2__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_2__2__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_2__2__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_2__2__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_2__2__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_2__2__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_1_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_0_ccff_tail));

	grid_io_right grid_io_right_3__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[24:31]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_2__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_2__1__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_2__1__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_2__1__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_2__1__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_2__1__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_2__1__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_2__1__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_0_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_1_ccff_tail));

	grid_io_bottom grid_io_bottom_2__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[32:39]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_2__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_2__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_2__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_2__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_2__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_2__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_2__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_2__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_0_ccff_tail));

	grid_io_bottom grid_io_bottom_1__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[40:47]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(ccff_head),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_1_ccff_tail));

	grid_io_left grid_io_left_0__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[48:55]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__0_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_0_ccff_tail));

	grid_io_left grid_io_left_0__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[56:63]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__1_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_1_ccff_tail));

	grid_clb grid_clb_1__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_1__1__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_clk_0_),
		.ccff_head(cby_1__1__0_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_0_ccff_tail));

	grid_clb grid_clb_1__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_1__2__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I_0_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_2_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.right_width_0_height_0_subtile_0__pin_I_3_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.right_width_0_height_0_subtile_0__pin_I_4_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_6_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.right_width_0_height_0_subtile_0__pin_I_7_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.right_width_0_height_0_subtile_0__pin_I_8_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_10_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.right_width_0_height_0_subtile_0__pin_I_11_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.right_width_0_height_0_subtile_0__pin_I_12_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_14_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.right_width_0_height_0_subtile_0__pin_I_15_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.right_width_0_height_0_subtile_0__pin_I_16_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_18_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.right_width_0_height_0_subtile_0__pin_I_19_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_clk_0_),
		.ccff_head(cby_1__2__0_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_0_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_3_),
		.right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_4_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_6_),
		.right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(ccff_tail));

	grid_memory grid_memory_2__1_ (
		.clk(clk),
		.right_width_0_height_0_subtile_0__pin_waddr_0_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_waddr_0_),
		.right_width_0_height_0_subtile_0__pin_waddr_1_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_waddr_1_),
		.right_width_0_height_0_subtile_0__pin_waddr_2_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.right_width_0_height_0_subtile_0__pin_waddr_3_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_waddr_3_),
		.right_width_0_height_0_subtile_0__pin_waddr_4_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_waddr_4_),
		.right_width_0_height_0_subtile_0__pin_raddr_0_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_raddr_0_),
		.right_width_0_height_0_subtile_0__pin_raddr_1_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.right_width_0_height_0_subtile_0__pin_raddr_2_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_raddr_2_),
		.right_width_0_height_0_subtile_0__pin_raddr_3_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_raddr_3_),
		.right_width_0_height_0_subtile_0__pin_raddr_4_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_raddr_4_),
		.right_width_0_height_0_subtile_0__pin_data_in_0_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.right_width_0_height_0_subtile_0__pin_data_in_1_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_data_in_1_),
		.right_width_0_height_0_subtile_0__pin_data_in_2_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_data_in_2_),
		.right_width_0_height_0_subtile_0__pin_data_in_3_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_data_in_3_),
		.right_width_0_height_0_subtile_0__pin_wen_0_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_5_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_5_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_6_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_6_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_7_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_7_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_8_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_8_),
		.bottom_width_0_height_0_subtile_0__pin_waddr_9_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_9_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_5_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_5_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_6_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_6_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_7_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_7_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_8_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_8_),
		.bottom_width_0_height_0_subtile_0__pin_raddr_9_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_9_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_4_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_4_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_5_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_5_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_6_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_6_),
		.bottom_width_0_height_0_subtile_0__pin_data_in_7_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_7_),
		.bottom_width_0_height_0_subtile_0__pin_ren_0_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ren_0_),
		.left_width_0_height_0_subtile_0__pin_clk_0_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_data_out_0_(grid_memory_0_right_width_0_height_0_subtile_0__pin_data_out_0_),
		.right_width_0_height_0_subtile_0__pin_data_out_1_(grid_memory_0_right_width_0_height_0_subtile_0__pin_data_out_1_),
		.right_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_0_right_width_0_height_0_subtile_0__pin_data_out_2_),
		.right_width_0_height_0_subtile_0__pin_data_out_3_(grid_memory_0_right_width_0_height_0_subtile_0__pin_data_out_3_),
		.bottom_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_0_bottom_width_0_height_0_subtile_0__pin_data_out_4_),
		.bottom_width_0_height_0_subtile_0__pin_data_out_5_(grid_memory_0_bottom_width_0_height_0_subtile_0__pin_data_out_5_),
		.bottom_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_0_bottom_width_0_height_0_subtile_0__pin_data_out_6_),
		.bottom_width_0_height_0_subtile_0__pin_data_out_7_(grid_memory_0_bottom_width_0_height_0_subtile_0__pin_data_out_7_));

	sb_0__0_ sb_0__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__0_chany_bottom_out[0:10]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__0__0_chanx_left_out[0:10]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_1_ccff_tail),
		.chany_top_out(sb_0__0__0_chany_top_out[0:10]),
		.chanx_right_out(sb_0__0__0_chanx_right_out[0:10]),
		.ccff_tail(sb_0__0__0_ccff_tail));

	sb_0__1_ sb_0__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__1_chany_bottom_out[0:10]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__0_chanx_left_out[0:10]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.chany_bottom_in(cby_0__1__0_chany_top_out[0:10]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_0__2__0_ccff_tail),
		.chany_top_out(sb_0__1__0_chany_top_out[0:10]),
		.chanx_right_out(sb_0__1__0_chanx_right_out[0:10]),
		.chany_bottom_out(sb_0__1__0_chany_bottom_out[0:10]),
		.ccff_tail(sb_0__1__0_ccff_tail));

	sb_0__2_ sb_0__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__2__0_chanx_left_out[0:10]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_0__1__1_chany_top_out[0:10]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_0_ccff_tail),
		.chanx_right_out(sb_0__2__0_chanx_right_out[0:10]),
		.chany_bottom_out(sb_0__2__0_chany_bottom_out[0:10]),
		.ccff_tail(sb_0__2__0_ccff_tail));

	sb_1__0_ sb_1__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__0_chany_bottom_out[0:10]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_right_in(cbx_2__0__0_chanx_left_out[0:10]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_0_bottom_width_0_height_0_subtile_0__pin_data_out_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_5_(grid_memory_0_bottom_width_0_height_0_subtile_0__pin_data_out_5_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_0_bottom_width_0_height_0_subtile_0__pin_data_out_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_7_(grid_memory_0_bottom_width_0_height_0_subtile_0__pin_data_out_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__0_chanx_right_out[0:10]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_0_ccff_tail),
		.chany_top_out(sb_1__0__0_chany_top_out[0:10]),
		.chanx_right_out(sb_1__0__0_chanx_right_out[0:10]),
		.chanx_left_out(sb_1__0__0_chanx_left_out[0:10]),
		.ccff_tail(sb_1__0__0_ccff_tail));

	sb_1__1_ sb_1__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__2__0_chany_bottom_out[0:10]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_),
		.chany_bottom_in(cby_1__1__0_chany_top_out[0:10]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(cbx_1__1__0_chanx_right_out[0:10]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_16_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_17_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_18_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_19_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_19_),
		.ccff_head(cby_2__2__0_ccff_tail),
		.chany_top_out(sb_1__1__0_chany_top_out[0:10]),
		.chany_bottom_out(sb_1__1__0_chany_bottom_out[0:10]),
		.chanx_left_out(sb_1__1__0_chanx_left_out[0:10]),
		.ccff_tail(sb_1__1__0_ccff_tail));

	sb_1__2_ sb_1__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__2__1_chanx_left_out[0:10]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_1__2__0_chany_top_out[0:10]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(cbx_1__2__0_chanx_right_out[0:10]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_1_ccff_tail),
		.chanx_right_out(sb_1__2__0_chanx_right_out[0:10]),
		.chany_bottom_out(sb_1__2__0_chany_bottom_out[0:10]),
		.chanx_left_out(sb_1__2__0_chanx_left_out[0:10]),
		.ccff_tail(sb_1__2__0_ccff_tail));

	sb_2__0_ sb_2__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_2__1__0_chany_bottom_out[0:10]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_0_(grid_memory_0_right_width_0_height_0_subtile_0__pin_data_out_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_1_(grid_memory_0_right_width_0_height_0_subtile_0__pin_data_out_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_0_right_width_0_height_0_subtile_0__pin_data_out_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_data_out_3_(grid_memory_0_right_width_0_height_0_subtile_0__pin_data_out_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_2__0__0_chanx_right_out[0:10]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_4_(grid_memory_0_bottom_width_0_height_0_subtile_0__pin_data_out_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_5_(grid_memory_0_bottom_width_0_height_0_subtile_0__pin_data_out_5_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_6_(grid_memory_0_bottom_width_0_height_0_subtile_0__pin_data_out_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_data_out_7_(grid_memory_0_bottom_width_0_height_0_subtile_0__pin_data_out_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_clb_0_ccff_tail),
		.chany_top_out(sb_2__0__0_chany_top_out[0:10]),
		.chanx_left_out(sb_2__0__0_chanx_left_out[0:10]),
		.ccff_tail(sb_2__0__0_ccff_tail));

	sb_2__1_ sb_2__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_2__2__0_chany_bottom_out[0:10]),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_2__1__0_chany_top_out[0:10]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_0_(grid_memory_0_right_width_0_height_0_subtile_0__pin_data_out_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_1_(grid_memory_0_right_width_0_height_0_subtile_0__pin_data_out_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_2_(grid_memory_0_right_width_0_height_0_subtile_0__pin_data_out_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_data_out_3_(grid_memory_0_right_width_0_height_0_subtile_0__pin_data_out_3_),
		.ccff_head(cby_2__1__0_ccff_tail),
		.chany_top_out(sb_2__1__0_chany_top_out[0:10]),
		.chany_bottom_out(sb_2__1__0_chany_bottom_out[0:10]),
		.ccff_tail(sb_2__1__0_ccff_tail));

	sb_2__2_ sb_2__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_2__2__0_chany_top_out[0:10]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__2__1_chanx_right_out[0:10]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_right_0_ccff_tail),
		.chany_bottom_out(sb_2__2__0_chany_bottom_out[0:10]),
		.chanx_left_out(sb_2__2__0_chanx_left_out[0:10]),
		.ccff_tail(sb_2__2__0_ccff_tail));

	cbx_1__0_ cbx_1__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__0__0_chanx_right_out[0:10]),
		.chanx_right_in(sb_1__0__0_chanx_left_out[0:10]),
		.ccff_head(sb_1__0__0_ccff_tail),
		.chanx_left_out(cbx_1__0__0_chanx_left_out[0:10]),
		.chanx_right_out(cbx_1__0__0_chanx_right_out[0:10]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__0_ccff_tail));

	cbx_1__1_ cbx_1__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__0_chanx_right_out[0:10]),
		.chanx_right_in(sb_1__1__0_chanx_left_out[0:10]),
		.ccff_head(sb_1__1__0_ccff_tail),
		.chanx_left_out(cbx_1__1__0_chanx_left_out[0:10]),
		.chanx_right_out(cbx_1__1__0_chanx_right_out[0:10]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_36_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_37_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_tail(cbx_1__1__0_ccff_tail));

	cbx_1__2_ cbx_1__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__2__0_chanx_right_out[0:10]),
		.chanx_right_in(sb_1__2__0_chanx_left_out[0:10]),
		.ccff_head(sb_1__2__0_ccff_tail),
		.chanx_left_out(cbx_1__2__0_chanx_left_out[0:10]),
		.chanx_right_out(cbx_1__2__0_chanx_right_out[0:10]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__2__0_ccff_tail));

	cbx_1__2_ cbx_2__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__2__0_chanx_right_out[0:10]),
		.chanx_right_in(sb_2__2__0_chanx_left_out[0:10]),
		.ccff_head(sb_2__2__0_ccff_tail),
		.chanx_left_out(cbx_1__2__1_chanx_left_out[0:10]),
		.chanx_right_out(cbx_1__2__1_chanx_right_out[0:10]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__2__1_ccff_tail));

	cbx_2__0_ cbx_2__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__0_chanx_right_out[0:10]),
		.chanx_right_in(sb_2__0__0_chanx_left_out[0:10]),
		.ccff_head(sb_2__0__0_ccff_tail),
		.chanx_left_out(cbx_2__0__0_chanx_left_out[0:10]),
		.chanx_right_out(cbx_2__0__0_chanx_right_out[0:10]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_5_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_6_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_7_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_8_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_8_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_9_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_waddr_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_5_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_6_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_7_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_8_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_8_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_9_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_raddr_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_4_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_5_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_6_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_7_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_data_in_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ren_0_(cbx_2__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ren_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_2__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_2__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_2__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_2__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_2__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_2__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_2__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_2__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_2__0__0_ccff_tail));

	cby_0__1_ cby_0__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__0__0_chany_top_out[0:10]),
		.chany_top_in(sb_0__1__0_chany_bottom_out[0:10]),
		.ccff_head(sb_0__0__0_ccff_tail),
		.chany_bottom_out(cby_0__1__0_chany_bottom_out[0:10]),
		.chany_top_out(cby_0__1__0_chany_top_out[0:10]),
		.right_grid_left_width_0_height_0_subtile_0__pin_clk_0_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_clk_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__0_ccff_tail));

	cby_0__1_ cby_0__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__0_chany_top_out[0:10]),
		.chany_top_in(sb_0__2__0_chany_bottom_out[0:10]),
		.ccff_head(sb_0__1__0_ccff_tail),
		.chany_bottom_out(cby_0__1__1_chany_bottom_out[0:10]),
		.chany_top_out(cby_0__1__1_chany_top_out[0:10]),
		.right_grid_left_width_0_height_0_subtile_0__pin_clk_0_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_clk_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__1_ccff_tail));

	cby_1__1_ cby_1__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__0_chany_top_out[0:10]),
		.chany_top_in(sb_1__1__0_chany_bottom_out[0:10]),
		.ccff_head(cbx_1__0__0_ccff_tail),
		.chany_bottom_out(cby_1__1__0_chany_bottom_out[0:10]),
		.chany_top_out(cby_1__1__0_chany_top_out[0:10]),
		.right_grid_left_width_0_height_0_subtile_0__pin_clk_0_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_clk_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_1__1__0_ccff_tail));

	cby_1__2_ cby_1__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__0_chany_top_out[0:10]),
		.chany_top_in(sb_1__2__0_chany_bottom_out[0:10]),
		.ccff_head(cbx_1__1__0_ccff_tail),
		.chany_bottom_out(cby_1__2__0_chany_bottom_out[0:10]),
		.chany_top_out(cby_1__2__0_chany_top_out[0:10]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_0_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_2_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_3_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_4_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_6_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_7_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_8_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_10_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_11_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_12_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_14_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_15_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_16_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_18_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_19_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_19_),
		.ccff_tail(cby_1__2__0_ccff_tail));

	cby_2__1_ cby_2__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_2__0__0_chany_top_out[0:10]),
		.chany_top_in(sb_2__1__0_chany_bottom_out[0:10]),
		.ccff_head(cbx_2__0__0_ccff_tail),
		.chany_bottom_out(cby_2__1__0_chany_bottom_out[0:10]),
		.chany_top_out(cby_2__1__0_chany_top_out[0:10]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_2__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_2__1__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_2__1__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_2__1__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_2__1__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_2__1__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_2__1__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_2__1__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_0_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_waddr_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_1_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_waddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_waddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_3_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_waddr_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_waddr_4_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_waddr_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_0_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_raddr_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_raddr_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_2_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_raddr_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_3_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_raddr_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_raddr_4_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_raddr_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_data_in_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_1_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_data_in_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_2_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_data_in_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_data_in_3_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_data_in_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_wen_0_(cby_2__1__0_left_grid_right_width_0_height_0_subtile_0__pin_wen_0_),
		.ccff_tail(cby_2__1__0_ccff_tail));

	cby_2__2_ cby_2__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_2__1__0_chany_top_out[0:10]),
		.chany_top_in(sb_2__2__0_chany_bottom_out[0:10]),
		.ccff_head(sb_2__1__0_ccff_tail),
		.chany_bottom_out(cby_2__2__0_chany_bottom_out[0:10]),
		.chany_top_out(cby_2__2__0_chany_top_out[0:10]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_2__2__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_2__2__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_2__2__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_2__2__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_2__2__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_2__2__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_2__2__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_2__2__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_2__2__0_ccff_tail));

endmodule
// ----- END Verilog module for fpga_top -----

//----- Default net type -----
`default_nettype none




